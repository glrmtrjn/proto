

library IEEE;
use IEEE.std_logic_1164.all;
use work.P_AES.all;
entity vezes is
	port(
		entrada : in std_logic_vector(7 downto 0);
		saida : out std_logic_vector(7 downto 0)
	);
end vezes;
----------------------
architecture dois of vezes is
	signal sinal : std_logic_vector(7 downto 0);  
begin
	sinal <= (others => entrada(7));
	saida <= (entrada(6 downto 0) &'0') xor (sinal and x"1b");

end dois;
----------------------
architecture tres of vezes is
	signal sinal : std_logic_vector(7 downto 0);
begin
	sinal <= (others => entrada(7));
	saida <= ((entrada(6 downto 0) &'0') xor entrada) xor (sinal and x"1b");

end tres;
----------------------
architecture nove of vezes is
begin
	
saida <=
	x"00" when entrada = x"00" else
	x"09" when entrada = x"01" else
	x"12" when entrada = x"02" else
	x"1b" when entrada = x"03" else
	x"24" when entrada = x"04" else
	x"2d" when entrada = x"05" else
	x"36" when entrada = x"06" else
	x"3f" when entrada = x"07" else
	x"48" when entrada = x"08" else
	x"41" when entrada = x"09" else
	x"5a" when entrada = x"0a" else
	x"53" when entrada = x"0b" else
	x"6c" when entrada = x"0c" else
	x"65" when entrada = x"0d" else
	x"7e" when entrada = x"0e" else
	x"77" when entrada = x"0f" else
	x"90" when entrada = x"10" else
	x"99" when entrada = x"11" else
	x"82" when entrada = x"12" else
	x"8b" when entrada = x"13" else
	x"b4" when entrada = x"14" else
	x"bd" when entrada = x"15" else
	x"a6" when entrada = x"16" else
	x"af" when entrada = x"17" else
	x"d8" when entrada = x"18" else
	x"d1" when entrada = x"19" else
	x"ca" when entrada = x"1a" else
	x"c3" when entrada = x"1b" else
	x"fc" when entrada = x"1c" else
	x"f5" when entrada = x"1d" else
	x"ee" when entrada = x"1e" else
	x"e7" when entrada = x"1f" else
	x"3b" when entrada = x"20" else
	x"32" when entrada = x"21" else
	x"29" when entrada = x"22" else
	x"20" when entrada = x"23" else
	x"1f" when entrada = x"24" else
	x"16" when entrada = x"25" else
	x"0d" when entrada = x"26" else
	x"04" when entrada = x"27" else
	x"73" when entrada = x"28" else
	x"7a" when entrada = x"29" else
	x"61" when entrada = x"2a" else
	x"68" when entrada = x"2b" else
	x"57" when entrada = x"2c" else
	x"5e" when entrada = x"2d" else
	x"45" when entrada = x"2e" else
	x"4c" when entrada = x"2f" else
	x"ab" when entrada = x"30" else
	x"a2" when entrada = x"31" else
	x"b9" when entrada = x"32" else
	x"b0" when entrada = x"33" else
	x"8f" when entrada = x"34" else
	x"86" when entrada = x"35" else
	x"9d" when entrada = x"36" else
	x"94" when entrada = x"37" else
	x"e3" when entrada = x"38" else
	x"ea" when entrada = x"39" else
	x"f1" when entrada = x"3a" else
	x"f8" when entrada = x"3b" else
	x"c7" when entrada = x"3c" else
	x"ce" when entrada = x"3d" else
	x"d5" when entrada = x"3e" else
	x"dc" when entrada = x"3f" else
	x"76" when entrada = x"40" else
	x"7f" when entrada = x"41" else
	x"64" when entrada = x"42" else
	x"6d" when entrada = x"43" else
	x"52" when entrada = x"44" else
	x"5b" when entrada = x"45" else
	x"40" when entrada = x"46" else
	x"49" when entrada = x"47" else
	x"3e" when entrada = x"48" else
	x"37" when entrada = x"49" else
	x"2c" when entrada = x"4a" else
	x"25" when entrada = x"4b" else
	x"1a" when entrada = x"4c" else
	x"13" when entrada = x"4d" else
	x"08" when entrada = x"4e" else
	x"01" when entrada = x"4f" else
	x"e6" when entrada = x"50" else
	x"ef" when entrada = x"51" else
	x"f4" when entrada = x"52" else
	x"fd" when entrada = x"53" else
	x"c2" when entrada = x"54" else
	x"cb" when entrada = x"55" else
	x"d0" when entrada = x"56" else
	x"d9" when entrada = x"57" else
	x"ae" when entrada = x"58" else
	x"a7" when entrada = x"59" else
	x"bc" when entrada = x"5a" else
	x"b5" when entrada = x"5b" else
	x"8a" when entrada = x"5c" else
	x"83" when entrada = x"5d" else
	x"98" when entrada = x"5e" else
	x"91" when entrada = x"5f" else
	x"4d" when entrada = x"60" else
	x"44" when entrada = x"61" else
	x"5f" when entrada = x"62" else
	x"56" when entrada = x"63" else
	x"69" when entrada = x"64" else
	x"60" when entrada = x"65" else
	x"7b" when entrada = x"66" else
	x"72" when entrada = x"67" else
	x"05" when entrada = x"68" else
	x"0c" when entrada = x"69" else
	x"17" when entrada = x"6a" else
	x"1e" when entrada = x"6b" else
	x"21" when entrada = x"6c" else
	x"28" when entrada = x"6d" else
	x"33" when entrada = x"6e" else
	x"3a" when entrada = x"6f" else
	x"dd" when entrada = x"70" else
	x"d4" when entrada = x"71" else
	x"cf" when entrada = x"72" else
	x"c6" when entrada = x"73" else
	x"f9" when entrada = x"74" else
	x"f0" when entrada = x"75" else
	x"eb" when entrada = x"76" else
	x"e2" when entrada = x"77" else
	x"95" when entrada = x"78" else
	x"9c" when entrada = x"79" else
	x"87" when entrada = x"7a" else
	x"8e" when entrada = x"7b" else
	x"b1" when entrada = x"7c" else
	x"b8" when entrada = x"7d" else
	x"a3" when entrada = x"7e" else
	x"aa" when entrada = x"7f" else
	x"ec" when entrada = x"80" else
	x"e5" when entrada = x"81" else
	x"fe" when entrada = x"82" else
	x"f7" when entrada = x"83" else
	x"c8" when entrada = x"84" else
	x"c1" when entrada = x"85" else
	x"da" when entrada = x"86" else
	x"d3" when entrada = x"87" else
	x"a4" when entrada = x"88" else
	x"ad" when entrada = x"89" else
	x"b6" when entrada = x"8a" else
	x"bf" when entrada = x"8b" else
	x"80" when entrada = x"8c" else
	x"89" when entrada = x"8d" else
	x"92" when entrada = x"8e" else
	x"9b" when entrada = x"8f" else
	x"7c" when entrada = x"90" else
	x"75" when entrada = x"91" else
	x"6e" when entrada = x"92" else
	x"67" when entrada = x"93" else
	x"58" when entrada = x"94" else
	x"51" when entrada = x"95" else
	x"4a" when entrada = x"96" else
	x"43" when entrada = x"97" else
	x"34" when entrada = x"98" else
	x"3d" when entrada = x"99" else
	x"26" when entrada = x"9a" else
	x"2f" when entrada = x"9b" else
	x"10" when entrada = x"9c" else
	x"19" when entrada = x"9d" else
	x"02" when entrada = x"9e" else
	x"0b" when entrada = x"9f" else
	x"d7" when entrada = x"a0" else
	x"de" when entrada = x"a1" else
	x"c5" when entrada = x"a2" else
	x"cc" when entrada = x"a3" else
	x"f3" when entrada = x"a4" else
	x"fa" when entrada = x"a5" else
	x"e1" when entrada = x"a6" else
	x"e8" when entrada = x"a7" else
	x"9f" when entrada = x"a8" else
	x"96" when entrada = x"a9" else
	x"8d" when entrada = x"aa" else
	x"84" when entrada = x"ab" else
	x"bb" when entrada = x"ac" else
	x"b2" when entrada = x"ad" else
	x"a9" when entrada = x"ae" else
	x"a0" when entrada = x"af" else
	x"47" when entrada = x"b0" else
	x"4e" when entrada = x"b1" else
	x"55" when entrada = x"b2" else
	x"5c" when entrada = x"b3" else
	x"63" when entrada = x"b4" else
	x"6a" when entrada = x"b5" else
	x"71" when entrada = x"b6" else
	x"78" when entrada = x"b7" else
	x"0f" when entrada = x"b8" else
	x"06" when entrada = x"b9" else
	x"1d" when entrada = x"ba" else
	x"14" when entrada = x"bb" else
	x"2b" when entrada = x"bc" else
	x"22" when entrada = x"bd" else
	x"39" when entrada = x"be" else
	x"30" when entrada = x"bf" else
	x"9a" when entrada = x"c0" else
	x"93" when entrada = x"c1" else
	x"88" when entrada = x"c2" else
	x"81" when entrada = x"c3" else
	x"be" when entrada = x"c4" else
	x"b7" when entrada = x"c5" else
	x"ac" when entrada = x"c6" else
	x"a5" when entrada = x"c7" else
	x"d2" when entrada = x"c8" else
	x"db" when entrada = x"c9" else
	x"c0" when entrada = x"ca" else
	x"c9" when entrada = x"cb" else
	x"f6" when entrada = x"cc" else
	x"ff" when entrada = x"cd" else
	x"e4" when entrada = x"ce" else
	x"ed" when entrada = x"cf" else
	x"0a" when entrada = x"d0" else
	x"03" when entrada = x"d1" else
	x"18" when entrada = x"d2" else
	x"11" when entrada = x"d3" else
	x"2e" when entrada = x"d4" else
	x"27" when entrada = x"d5" else
	x"3c" when entrada = x"d6" else
	x"35" when entrada = x"d7" else
	x"42" when entrada = x"d8" else
	x"4b" when entrada = x"d9" else
	x"50" when entrada = x"da" else
	x"59" when entrada = x"db" else
	x"66" when entrada = x"dc" else
	x"6f" when entrada = x"dd" else
	x"74" when entrada = x"de" else
	x"7d" when entrada = x"df" else
	x"a1" when entrada = x"e0" else
	x"a8" when entrada = x"e1" else
	x"b3" when entrada = x"e2" else
	x"ba" when entrada = x"e3" else
	x"85" when entrada = x"e4" else
	x"8c" when entrada = x"e5" else
	x"97" when entrada = x"e6" else
	x"9e" when entrada = x"e7" else
	x"e9" when entrada = x"e8" else
	x"e0" when entrada = x"e9" else
	x"fb" when entrada = x"ea" else
	x"f2" when entrada = x"eb" else
	x"cd" when entrada = x"ec" else
	x"c4" when entrada = x"ed" else
	x"df" when entrada = x"ee" else
	x"d6" when entrada = x"ef" else
	x"31" when entrada = x"f0" else
	x"38" when entrada = x"f1" else
	x"23" when entrada = x"f2" else
	x"2a" when entrada = x"f3" else
	x"15" when entrada = x"f4" else
	x"1c" when entrada = x"f5" else
	x"07" when entrada = x"f6" else
	x"0e" when entrada = x"f7" else
	x"79" when entrada = x"f8" else
	x"70" when entrada = x"f9" else
	x"6b" when entrada = x"fa" else
	x"62" when entrada = x"fb" else
	x"5d" when entrada = x"fc" else
	x"54" when entrada = x"fd" else
	x"4f" when entrada = x"fe" else
	x"46" when entrada = x"ff";

end nove;
----------------------
architecture onze of vezes is
begin
saida <=
	x"00" when entrada = x"00" else
	x"0b" when entrada = x"01" else
	x"16" when entrada = x"02" else
	x"1d" when entrada = x"03" else
	x"2c" when entrada = x"04" else
	x"27" when entrada = x"05" else
	x"3a" when entrada = x"06" else
	x"31" when entrada = x"07" else
	x"58" when entrada = x"08" else
	x"53" when entrada = x"09" else
	x"4e" when entrada = x"0a" else
	x"45" when entrada = x"0b" else
	x"74" when entrada = x"0c" else
	x"7f" when entrada = x"0d" else
	x"62" when entrada = x"0e" else
	x"69" when entrada = x"0f" else
	x"b0" when entrada = x"10" else
	x"bb" when entrada = x"11" else
	x"a6" when entrada = x"12" else
	x"ad" when entrada = x"13" else
	x"9c" when entrada = x"14" else
	x"97" when entrada = x"15" else
	x"8a" when entrada = x"16" else
	x"81" when entrada = x"17" else
	x"e8" when entrada = x"18" else
	x"e3" when entrada = x"19" else
	x"fe" when entrada = x"1a" else
	x"f5" when entrada = x"1b" else
	x"c4" when entrada = x"1c" else
	x"cf" when entrada = x"1d" else
	x"d2" when entrada = x"1e" else
	x"d9" when entrada = x"1f" else
	x"7b" when entrada = x"20" else
	x"70" when entrada = x"21" else
	x"6d" when entrada = x"22" else
	x"66" when entrada = x"23" else
	x"57" when entrada = x"24" else
	x"5c" when entrada = x"25" else
	x"41" when entrada = x"26" else
	x"4a" when entrada = x"27" else
	x"23" when entrada = x"28" else
	x"28" when entrada = x"29" else
	x"35" when entrada = x"2a" else
	x"3e" when entrada = x"2b" else
	x"0f" when entrada = x"2c" else
	x"04" when entrada = x"2d" else
	x"19" when entrada = x"2e" else
	x"12" when entrada = x"2f" else
	x"cb" when entrada = x"30" else
	x"c0" when entrada = x"31" else
	x"dd" when entrada = x"32" else
	x"d6" when entrada = x"33" else
	x"e7" when entrada = x"34" else
	x"ec" when entrada = x"35" else
	x"f1" when entrada = x"36" else
	x"fa" when entrada = x"37" else
	x"93" when entrada = x"38" else
	x"98" when entrada = x"39" else
	x"85" when entrada = x"3a" else
	x"8e" when entrada = x"3b" else
	x"bf" when entrada = x"3c" else
	x"b4" when entrada = x"3d" else
	x"a9" when entrada = x"3e" else
	x"a2" when entrada = x"3f" else
	x"f6" when entrada = x"40" else
	x"fd" when entrada = x"41" else
	x"e0" when entrada = x"42" else
	x"eb" when entrada = x"43" else
	x"da" when entrada = x"44" else
	x"d1" when entrada = x"45" else
	x"cc" when entrada = x"46" else
	x"c7" when entrada = x"47" else
	x"ae" when entrada = x"48" else
	x"a5" when entrada = x"49" else
	x"b8" when entrada = x"4a" else
	x"b3" when entrada = x"4b" else
	x"82" when entrada = x"4c" else
	x"89" when entrada = x"4d" else
	x"94" when entrada = x"4e" else
	x"9f" when entrada = x"4f" else
	x"46" when entrada = x"50" else
	x"4d" when entrada = x"51" else
	x"50" when entrada = x"52" else
	x"5b" when entrada = x"53" else
	x"6a" when entrada = x"54" else
	x"61" when entrada = x"55" else
	x"7c" when entrada = x"56" else
	x"77" when entrada = x"57" else
	x"1e" when entrada = x"58" else
	x"15" when entrada = x"59" else
	x"08" when entrada = x"5a" else
	x"03" when entrada = x"5b" else
	x"32" when entrada = x"5c" else
	x"39" when entrada = x"5d" else
	x"24" when entrada = x"5e" else
	x"2f" when entrada = x"5f" else
	x"8d" when entrada = x"60" else
	x"86" when entrada = x"61" else
	x"9b" when entrada = x"62" else
	x"90" when entrada = x"63" else
	x"a1" when entrada = x"64" else
	x"aa" when entrada = x"65" else
	x"b7" when entrada = x"66" else
	x"bc" when entrada = x"67" else
	x"d5" when entrada = x"68" else
	x"de" when entrada = x"69" else
	x"c3" when entrada = x"6a" else
	x"c8" when entrada = x"6b" else
	x"f9" when entrada = x"6c" else
	x"f2" when entrada = x"6d" else
	x"ef" when entrada = x"6e" else
	x"e4" when entrada = x"6f" else
	x"3d" when entrada = x"70" else
	x"36" when entrada = x"71" else
	x"2b" when entrada = x"72" else
	x"20" when entrada = x"73" else
	x"11" when entrada = x"74" else
	x"1a" when entrada = x"75" else
	x"07" when entrada = x"76" else
	x"0c" when entrada = x"77" else
	x"65" when entrada = x"78" else
	x"6e" when entrada = x"79" else
	x"73" when entrada = x"7a" else
	x"78" when entrada = x"7b" else
	x"49" when entrada = x"7c" else
	x"42" when entrada = x"7d" else
	x"5f" when entrada = x"7e" else
	x"54" when entrada = x"7f" else
	x"f7" when entrada = x"80" else
	x"fc" when entrada = x"81" else
	x"e1" when entrada = x"82" else
	x"ea" when entrada = x"83" else
	x"db" when entrada = x"84" else
	x"d0" when entrada = x"85" else
	x"cd" when entrada = x"86" else
	x"c6" when entrada = x"87" else
	x"af" when entrada = x"88" else
	x"a4" when entrada = x"89" else
	x"b9" when entrada = x"8a" else
	x"b2" when entrada = x"8b" else
	x"83" when entrada = x"8c" else
	x"88" when entrada = x"8d" else
	x"95" when entrada = x"8e" else
	x"9e" when entrada = x"8f" else
	x"47" when entrada = x"90" else
	x"4c" when entrada = x"91" else
	x"51" when entrada = x"92" else
	x"5a" when entrada = x"93" else
	x"6b" when entrada = x"94" else
	x"60" when entrada = x"95" else
	x"7d" when entrada = x"96" else
	x"76" when entrada = x"97" else
	x"1f" when entrada = x"98" else
	x"14" when entrada = x"99" else
	x"09" when entrada = x"9a" else
	x"02" when entrada = x"9b" else
	x"33" when entrada = x"9c" else
	x"38" when entrada = x"9d" else
	x"25" when entrada = x"9e" else
	x"2e" when entrada = x"9f" else
	x"8c" when entrada = x"a0" else
	x"87" when entrada = x"a1" else
	x"9a" when entrada = x"a2" else
	x"91" when entrada = x"a3" else
	x"a0" when entrada = x"a4" else
	x"ab" when entrada = x"a5" else
	x"b6" when entrada = x"a6" else
	x"bd" when entrada = x"a7" else
	x"d4" when entrada = x"a8" else
	x"df" when entrada = x"a9" else
	x"c2" when entrada = x"aa" else
	x"c9" when entrada = x"ab" else
	x"f8" when entrada = x"ac" else
	x"f3" when entrada = x"ad" else
	x"ee" when entrada = x"ae" else
	x"e5" when entrada = x"af" else
	x"3c" when entrada = x"b0" else
	x"37" when entrada = x"b1" else
	x"2a" when entrada = x"b2" else
	x"21" when entrada = x"b3" else
	x"10" when entrada = x"b4" else
	x"1b" when entrada = x"b5" else
	x"06" when entrada = x"b6" else
	x"0d" when entrada = x"b7" else
	x"64" when entrada = x"b8" else
	x"6f" when entrada = x"b9" else
	x"72" when entrada = x"ba" else
	x"79" when entrada = x"bb" else
	x"48" when entrada = x"bc" else
	x"43" when entrada = x"bd" else
	x"5e" when entrada = x"be" else
	x"55" when entrada = x"bf" else
	x"01" when entrada = x"c0" else
	x"0a" when entrada = x"c1" else
	x"17" when entrada = x"c2" else
	x"1c" when entrada = x"c3" else
	x"2d" when entrada = x"c4" else
	x"26" when entrada = x"c5" else
	x"3b" when entrada = x"c6" else
	x"30" when entrada = x"c7" else
	x"59" when entrada = x"c8" else
	x"52" when entrada = x"c9" else
	x"4f" when entrada = x"ca" else
	x"44" when entrada = x"cb" else
	x"75" when entrada = x"cc" else
	x"7e" when entrada = x"cd" else
	x"63" when entrada = x"ce" else
	x"68" when entrada = x"cf" else
	x"b1" when entrada = x"d0" else
	x"ba" when entrada = x"d1" else
	x"a7" when entrada = x"d2" else
	x"ac" when entrada = x"d3" else
	x"9d" when entrada = x"d4" else
	x"96" when entrada = x"d5" else
	x"8b" when entrada = x"d6" else
	x"80" when entrada = x"d7" else
	x"e9" when entrada = x"d8" else
	x"e2" when entrada = x"d9" else
	x"ff" when entrada = x"da" else
	x"f4" when entrada = x"db" else
	x"c5" when entrada = x"dc" else
	x"ce" when entrada = x"dd" else
	x"d3" when entrada = x"de" else
	x"d8" when entrada = x"df" else
	x"7a" when entrada = x"e0" else
	x"71" when entrada = x"e1" else
	x"6c" when entrada = x"e2" else
	x"67" when entrada = x"e3" else
	x"56" when entrada = x"e4" else
	x"5d" when entrada = x"e5" else
	x"40" when entrada = x"e6" else
	x"4b" when entrada = x"e7" else
	x"22" when entrada = x"e8" else
	x"29" when entrada = x"e9" else
	x"34" when entrada = x"ea" else
	x"3f" when entrada = x"eb" else
	x"0e" when entrada = x"ec" else
	x"05" when entrada = x"ed" else
	x"18" when entrada = x"ee" else
	x"13" when entrada = x"ef" else
	x"ca" when entrada = x"f0" else
	x"c1" when entrada = x"f1" else
	x"dc" when entrada = x"f2" else
	x"d7" when entrada = x"f3" else
	x"e6" when entrada = x"f4" else
	x"ed" when entrada = x"f5" else
	x"f0" when entrada = x"f6" else
	x"fb" when entrada = x"f7" else
	x"92" when entrada = x"f8" else
	x"99" when entrada = x"f9" else
	x"84" when entrada = x"fa" else
	x"8f" when entrada = x"fb" else
	x"be" when entrada = x"fc" else
	x"b5" when entrada = x"fd" else
	x"a8" when entrada = x"fe" else
	x"a3" when entrada = x"ff";	
end onze;
----------------------
architecture treze of vezes is
begin

saida <=
	x"00" when entrada = x"00" else
	x"0d" when entrada = x"01" else
	x"1a" when entrada = x"02" else
	x"17" when entrada = x"03" else
	x"34" when entrada = x"04" else
	x"39" when entrada = x"05" else
	x"2e" when entrada = x"06" else
	x"23" when entrada = x"07" else
	x"68" when entrada = x"08" else
	x"65" when entrada = x"09" else
	x"72" when entrada = x"0a" else
	x"7f" when entrada = x"0b" else
	x"5c" when entrada = x"0c" else
	x"51" when entrada = x"0d" else
	x"46" when entrada = x"0e" else
	x"4b" when entrada = x"0f" else
	x"d0" when entrada = x"10" else
	x"dd" when entrada = x"11" else
	x"ca" when entrada = x"12" else
	x"c7" when entrada = x"13" else
	x"e4" when entrada = x"14" else
	x"e9" when entrada = x"15" else
	x"fe" when entrada = x"16" else
	x"f3" when entrada = x"17" else
	x"b8" when entrada = x"18" else
	x"b5" when entrada = x"19" else
	x"a2" when entrada = x"1a" else
	x"af" when entrada = x"1b" else
	x"8c" when entrada = x"1c" else
	x"81" when entrada = x"1d" else
	x"96" when entrada = x"1e" else
	x"9b" when entrada = x"1f" else
	x"bb" when entrada = x"20" else
	x"b6" when entrada = x"21" else
	x"a1" when entrada = x"22" else
	x"ac" when entrada = x"23" else
	x"8f" when entrada = x"24" else
	x"82" when entrada = x"25" else
	x"95" when entrada = x"26" else
	x"98" when entrada = x"27" else
	x"d3" when entrada = x"28" else
	x"de" when entrada = x"29" else
	x"c9" when entrada = x"2a" else
	x"c4" when entrada = x"2b" else
	x"e7" when entrada = x"2c" else
	x"ea" when entrada = x"2d" else
	x"fd" when entrada = x"2e" else
	x"f0" when entrada = x"2f" else
	x"6b" when entrada = x"30" else
	x"66" when entrada = x"31" else
	x"71" when entrada = x"32" else
	x"7c" when entrada = x"33" else
	x"5f" when entrada = x"34" else
	x"52" when entrada = x"35" else
	x"45" when entrada = x"36" else
	x"48" when entrada = x"37" else
	x"03" when entrada = x"38" else
	x"0e" when entrada = x"39" else
	x"19" when entrada = x"3a" else
	x"14" when entrada = x"3b" else
	x"37" when entrada = x"3c" else
	x"3a" when entrada = x"3d" else
	x"2d" when entrada = x"3e" else
	x"20" when entrada = x"3f" else
	x"6d" when entrada = x"40" else
	x"60" when entrada = x"41" else
	x"77" when entrada = x"42" else
	x"7a" when entrada = x"43" else
	x"59" when entrada = x"44" else
	x"54" when entrada = x"45" else
	x"43" when entrada = x"46" else
	x"4e" when entrada = x"47" else
	x"05" when entrada = x"48" else
	x"08" when entrada = x"49" else
	x"1f" when entrada = x"4a" else
	x"12" when entrada = x"4b" else
	x"31" when entrada = x"4c" else
	x"3c" when entrada = x"4d" else
	x"2b" when entrada = x"4e" else
	x"26" when entrada = x"4f" else
	x"bd" when entrada = x"50" else
	x"b0" when entrada = x"51" else
	x"a7" when entrada = x"52" else
	x"aa" when entrada = x"53" else
	x"89" when entrada = x"54" else
	x"84" when entrada = x"55" else
	x"93" when entrada = x"56" else
	x"9e" when entrada = x"57" else
	x"d5" when entrada = x"58" else
	x"d8" when entrada = x"59" else
	x"cf" when entrada = x"5a" else
	x"c2" when entrada = x"5b" else
	x"e1" when entrada = x"5c" else
	x"ec" when entrada = x"5d" else
	x"fb" when entrada = x"5e" else
	x"f6" when entrada = x"5f" else
	x"d6" when entrada = x"60" else
	x"db" when entrada = x"61" else
	x"cc" when entrada = x"62" else
	x"c1" when entrada = x"63" else
	x"e2" when entrada = x"64" else
	x"ef" when entrada = x"65" else
	x"f8" when entrada = x"66" else
	x"f5" when entrada = x"67" else
	x"be" when entrada = x"68" else
	x"b3" when entrada = x"69" else
	x"a4" when entrada = x"6a" else
	x"a9" when entrada = x"6b" else
	x"8a" when entrada = x"6c" else
	x"87" when entrada = x"6d" else
	x"90" when entrada = x"6e" else
	x"9d" when entrada = x"6f" else
	x"06" when entrada = x"70" else
	x"0b" when entrada = x"71" else
	x"1c" when entrada = x"72" else
	x"11" when entrada = x"73" else
	x"32" when entrada = x"74" else
	x"3f" when entrada = x"75" else
	x"28" when entrada = x"76" else
	x"25" when entrada = x"77" else
	x"6e" when entrada = x"78" else
	x"63" when entrada = x"79" else
	x"74" when entrada = x"7a" else
	x"79" when entrada = x"7b" else
	x"5a" when entrada = x"7c" else
	x"57" when entrada = x"7d" else
	x"40" when entrada = x"7e" else
	x"4d" when entrada = x"7f" else
	x"da" when entrada = x"80" else
	x"d7" when entrada = x"81" else
	x"c0" when entrada = x"82" else
	x"cd" when entrada = x"83" else
	x"ee" when entrada = x"84" else
	x"e3" when entrada = x"85" else
	x"f4" when entrada = x"86" else
	x"f9" when entrada = x"87" else
	x"b2" when entrada = x"88" else
	x"bf" when entrada = x"89" else
	x"a8" when entrada = x"8a" else
	x"a5" when entrada = x"8b" else
	x"86" when entrada = x"8c" else
	x"8b" when entrada = x"8d" else
	x"9c" when entrada = x"8e" else
	x"91" when entrada = x"8f" else
	x"0a" when entrada = x"90" else
	x"07" when entrada = x"91" else
	x"10" when entrada = x"92" else
	x"1d" when entrada = x"93" else
	x"3e" when entrada = x"94" else
	x"33" when entrada = x"95" else
	x"24" when entrada = x"96" else
	x"29" when entrada = x"97" else
	x"62" when entrada = x"98" else
	x"6f" when entrada = x"99" else
	x"78" when entrada = x"9a" else
	x"75" when entrada = x"9b" else
	x"56" when entrada = x"9c" else
	x"5b" when entrada = x"9d" else
	x"4c" when entrada = x"9e" else
	x"41" when entrada = x"9f" else
	x"61" when entrada = x"a0" else
	x"6c" when entrada = x"a1" else
	x"7b" when entrada = x"a2" else
	x"76" when entrada = x"a3" else
	x"55" when entrada = x"a4" else
	x"58" when entrada = x"a5" else
	x"4f" when entrada = x"a6" else
	x"42" when entrada = x"a7" else
	x"09" when entrada = x"a8" else
	x"04" when entrada = x"a9" else
	x"13" when entrada = x"aa" else
	x"1e" when entrada = x"ab" else
	x"3d" when entrada = x"ac" else
	x"30" when entrada = x"ad" else
	x"27" when entrada = x"ae" else
	x"2a" when entrada = x"af" else
	x"b1" when entrada = x"b0" else
	x"bc" when entrada = x"b1" else
	x"ab" when entrada = x"b2" else
	x"a6" when entrada = x"b3" else
	x"85" when entrada = x"b4" else
	x"88" when entrada = x"b5" else
	x"9f" when entrada = x"b6" else
	x"92" when entrada = x"b7" else
	x"d9" when entrada = x"b8" else
	x"d4" when entrada = x"b9" else
	x"c3" when entrada = x"ba" else
	x"ce" when entrada = x"bb" else
	x"ed" when entrada = x"bc" else
	x"e0" when entrada = x"bd" else
	x"f7" when entrada = x"be" else
	x"fa" when entrada = x"bf" else
	x"b7" when entrada = x"c0" else
	x"ba" when entrada = x"c1" else
	x"ad" when entrada = x"c2" else
	x"a0" when entrada = x"c3" else
	x"83" when entrada = x"c4" else
	x"8e" when entrada = x"c5" else
	x"99" when entrada = x"c6" else
	x"94" when entrada = x"c7" else
	x"df" when entrada = x"c8" else
	x"d2" when entrada = x"c9" else
	x"c5" when entrada = x"ca" else
	x"c8" when entrada = x"cb" else
	x"eb" when entrada = x"cc" else
	x"e6" when entrada = x"cd" else
	x"f1" when entrada = x"ce" else
	x"fc" when entrada = x"cf" else
	x"67" when entrada = x"d0" else
	x"6a" when entrada = x"d1" else
	x"7d" when entrada = x"d2" else
	x"70" when entrada = x"d3" else
	x"53" when entrada = x"d4" else
	x"5e" when entrada = x"d5" else
	x"49" when entrada = x"d6" else
	x"44" when entrada = x"d7" else
	x"0f" when entrada = x"d8" else
	x"02" when entrada = x"d9" else
	x"15" when entrada = x"da" else
	x"18" when entrada = x"db" else
	x"3b" when entrada = x"dc" else
	x"36" when entrada = x"dd" else
	x"21" when entrada = x"de" else
	x"2c" when entrada = x"df" else
	x"0c" when entrada = x"e0" else
	x"01" when entrada = x"e1" else
	x"16" when entrada = x"e2" else
	x"1b" when entrada = x"e3" else
	x"38" when entrada = x"e4" else
	x"35" when entrada = x"e5" else
	x"22" when entrada = x"e6" else
	x"2f" when entrada = x"e7" else
	x"64" when entrada = x"e8" else
	x"69" when entrada = x"e9" else
	x"7e" when entrada = x"ea" else
	x"73" when entrada = x"eb" else
	x"50" when entrada = x"ec" else
	x"5d" when entrada = x"ed" else
	x"4a" when entrada = x"ee" else
	x"47" when entrada = x"ef" else
	x"dc" when entrada = x"f0" else
	x"d1" when entrada = x"f1" else
	x"c6" when entrada = x"f2" else
	x"cb" when entrada = x"f3" else
	x"e8" when entrada = x"f4" else
	x"e5" when entrada = x"f5" else
	x"f2" when entrada = x"f6" else
	x"ff" when entrada = x"f7" else
	x"b4" when entrada = x"f8" else
	x"b9" when entrada = x"f9" else
	x"ae" when entrada = x"fa" else
	x"a3" when entrada = x"fb" else
	x"80" when entrada = x"fc" else
	x"8d" when entrada = x"fd" else
	x"9a" when entrada = x"fe" else
	x"97" when entrada = x"ff";
	
end treze;
----------------------
architecture catorze of vezes is
begin
saida <=
	x"00" when entrada = x"00" else
	x"0e" when entrada = x"01" else
	x"1c" when entrada = x"02" else
	x"12" when entrada = x"03" else
	x"38" when entrada = x"04" else
	x"36" when entrada = x"05" else
	x"24" when entrada = x"06" else
	x"2a" when entrada = x"07" else
	x"70" when entrada = x"08" else
	x"7e" when entrada = x"09" else
	x"6c" when entrada = x"0a" else
	x"62" when entrada = x"0b" else
	x"48" when entrada = x"0c" else
	x"46" when entrada = x"0d" else
	x"54" when entrada = x"0e" else
	x"5a" when entrada = x"0f" else
	x"e0" when entrada = x"10" else
	x"ee" when entrada = x"11" else
	x"fc" when entrada = x"12" else
	x"f2" when entrada = x"13" else
	x"d8" when entrada = x"14" else
	x"d6" when entrada = x"15" else
	x"c4" when entrada = x"16" else
	x"ca" when entrada = x"17" else
	x"90" when entrada = x"18" else
	x"9e" when entrada = x"19" else
	x"8c" when entrada = x"1a" else
	x"82" when entrada = x"1b" else
	x"a8" when entrada = x"1c" else
	x"a6" when entrada = x"1d" else
	x"b4" when entrada = x"1e" else
	x"ba" when entrada = x"1f" else
	x"db" when entrada = x"20" else
	x"d5" when entrada = x"21" else
	x"c7" when entrada = x"22" else
	x"c9" when entrada = x"23" else
	x"e3" when entrada = x"24" else
	x"ed" when entrada = x"25" else
	x"ff" when entrada = x"26" else
	x"f1" when entrada = x"27" else
	x"ab" when entrada = x"28" else
	x"a5" when entrada = x"29" else
	x"b7" when entrada = x"2a" else
	x"b9" when entrada = x"2b" else
	x"93" when entrada = x"2c" else
	x"9d" when entrada = x"2d" else
	x"8f" when entrada = x"2e" else
	x"81" when entrada = x"2f" else
	x"3b" when entrada = x"30" else
	x"35" when entrada = x"31" else
	x"27" when entrada = x"32" else
	x"29" when entrada = x"33" else
	x"03" when entrada = x"34" else
	x"0d" when entrada = x"35" else
	x"1f" when entrada = x"36" else
	x"11" when entrada = x"37" else
	x"4b" when entrada = x"38" else
	x"45" when entrada = x"39" else
	x"57" when entrada = x"3a" else
	x"59" when entrada = x"3b" else
	x"73" when entrada = x"3c" else
	x"7d" when entrada = x"3d" else
	x"6f" when entrada = x"3e" else
	x"61" when entrada = x"3f" else
	x"ad" when entrada = x"40" else
	x"a3" when entrada = x"41" else
	x"b1" when entrada = x"42" else
	x"bf" when entrada = x"43" else
	x"95" when entrada = x"44" else
	x"9b" when entrada = x"45" else
	x"89" when entrada = x"46" else
	x"87" when entrada = x"47" else
	x"dd" when entrada = x"48" else
	x"d3" when entrada = x"49" else
	x"c1" when entrada = x"4a" else
	x"cf" when entrada = x"4b" else
	x"e5" when entrada = x"4c" else
	x"eb" when entrada = x"4d" else
	x"f9" when entrada = x"4e" else
	x"f7" when entrada = x"4f" else
	x"4d" when entrada = x"50" else
	x"43" when entrada = x"51" else
	x"51" when entrada = x"52" else
	x"5f" when entrada = x"53" else
	x"75" when entrada = x"54" else
	x"7b" when entrada = x"55" else
	x"69" when entrada = x"56" else
	x"67" when entrada = x"57" else
	x"3d" when entrada = x"58" else
	x"33" when entrada = x"59" else
	x"21" when entrada = x"5a" else
	x"2f" when entrada = x"5b" else
	x"05" when entrada = x"5c" else
	x"0b" when entrada = x"5d" else
	x"19" when entrada = x"5e" else
	x"17" when entrada = x"5f" else
	x"76" when entrada = x"60" else
	x"78" when entrada = x"61" else
	x"6a" when entrada = x"62" else
	x"64" when entrada = x"63" else
	x"4e" when entrada = x"64" else
	x"40" when entrada = x"65" else
	x"52" when entrada = x"66" else
	x"5c" when entrada = x"67" else
	x"06" when entrada = x"68" else
	x"08" when entrada = x"69" else
	x"1a" when entrada = x"6a" else
	x"14" when entrada = x"6b" else
	x"3e" when entrada = x"6c" else
	x"30" when entrada = x"6d" else
	x"22" when entrada = x"6e" else
	x"2c" when entrada = x"6f" else
	x"96" when entrada = x"70" else
	x"98" when entrada = x"71" else
	x"8a" when entrada = x"72" else
	x"84" when entrada = x"73" else
	x"ae" when entrada = x"74" else
	x"a0" when entrada = x"75" else
	x"b2" when entrada = x"76" else
	x"bc" when entrada = x"77" else
	x"e6" when entrada = x"78" else
	x"e8" when entrada = x"79" else
	x"fa" when entrada = x"7a" else
	x"f4" when entrada = x"7b" else
	x"de" when entrada = x"7c" else
	x"d0" when entrada = x"7d" else
	x"c2" when entrada = x"7e" else
	x"cc" when entrada = x"7f" else
	x"41" when entrada = x"80" else
	x"4f" when entrada = x"81" else
	x"5d" when entrada = x"82" else
	x"53" when entrada = x"83" else
	x"79" when entrada = x"84" else
	x"77" when entrada = x"85" else
	x"65" when entrada = x"86" else
	x"6b" when entrada = x"87" else
	x"31" when entrada = x"88" else
	x"3f" when entrada = x"89" else
	x"2d" when entrada = x"8a" else
	x"23" when entrada = x"8b" else
	x"09" when entrada = x"8c" else
	x"07" when entrada = x"8d" else
	x"15" when entrada = x"8e" else
	x"1b" when entrada = x"8f" else
	x"a1" when entrada = x"90" else
	x"af" when entrada = x"91" else
	x"bd" when entrada = x"92" else
	x"b3" when entrada = x"93" else
	x"99" when entrada = x"94" else
	x"97" when entrada = x"95" else
	x"85" when entrada = x"96" else
	x"8b" when entrada = x"97" else
	x"d1" when entrada = x"98" else
	x"df" when entrada = x"99" else
	x"cd" when entrada = x"9a" else
	x"c3" when entrada = x"9b" else
	x"e9" when entrada = x"9c" else
	x"e7" when entrada = x"9d" else
	x"f5" when entrada = x"9e" else
	x"fb" when entrada = x"9f" else
	x"9a" when entrada = x"a0" else
	x"94" when entrada = x"a1" else
	x"86" when entrada = x"a2" else
	x"88" when entrada = x"a3" else
	x"a2" when entrada = x"a4" else
	x"ac" when entrada = x"a5" else
	x"be" when entrada = x"a6" else
	x"b0" when entrada = x"a7" else
	x"ea" when entrada = x"a8" else
	x"e4" when entrada = x"a9" else
	x"f6" when entrada = x"aa" else
	x"f8" when entrada = x"ab" else
	x"d2" when entrada = x"ac" else
	x"dc" when entrada = x"ad" else
	x"ce" when entrada = x"ae" else
	x"c0" when entrada = x"af" else
	x"7a" when entrada = x"b0" else
	x"74" when entrada = x"b1" else
	x"66" when entrada = x"b2" else
	x"68" when entrada = x"b3" else
	x"42" when entrada = x"b4" else
	x"4c" when entrada = x"b5" else
	x"5e" when entrada = x"b6" else
	x"50" when entrada = x"b7" else
	x"0a" when entrada = x"b8" else
	x"04" when entrada = x"b9" else
	x"16" when entrada = x"ba" else
	x"18" when entrada = x"bb" else
	x"32" when entrada = x"bc" else
	x"3c" when entrada = x"bd" else
	x"2e" when entrada = x"be" else
	x"20" when entrada = x"bf" else
	x"ec" when entrada = x"c0" else
	x"e2" when entrada = x"c1" else
	x"f0" when entrada = x"c2" else
	x"fe" when entrada = x"c3" else
	x"d4" when entrada = x"c4" else
	x"da" when entrada = x"c5" else
	x"c8" when entrada = x"c6" else
	x"c6" when entrada = x"c7" else
	x"9c" when entrada = x"c8" else
	x"92" when entrada = x"c9" else
	x"80" when entrada = x"ca" else
	x"8e" when entrada = x"cb" else
	x"a4" when entrada = x"cc" else
	x"aa" when entrada = x"cd" else
	x"b8" when entrada = x"ce" else
	x"b6" when entrada = x"cf" else
	x"0c" when entrada = x"d0" else
	x"02" when entrada = x"d1" else
	x"10" when entrada = x"d2" else
	x"1e" when entrada = x"d3" else
	x"34" when entrada = x"d4" else
	x"3a" when entrada = x"d5" else
	x"28" when entrada = x"d6" else
	x"26" when entrada = x"d7" else
	x"7c" when entrada = x"d8" else
	x"72" when entrada = x"d9" else
	x"60" when entrada = x"da" else
	x"6e" when entrada = x"db" else
	x"44" when entrada = x"dc" else
	x"4a" when entrada = x"dd" else
	x"58" when entrada = x"de" else
	x"56" when entrada = x"df" else
	x"37" when entrada = x"e0" else
	x"39" when entrada = x"e1" else
	x"2b" when entrada = x"e2" else
	x"25" when entrada = x"e3" else
	x"0f" when entrada = x"e4" else
	x"01" when entrada = x"e5" else
	x"13" when entrada = x"e6" else
	x"1d" when entrada = x"e7" else
	x"47" when entrada = x"e8" else
	x"49" when entrada = x"e9" else
	x"5b" when entrada = x"ea" else
	x"55" when entrada = x"eb" else
	x"7f" when entrada = x"ec" else
	x"71" when entrada = x"ed" else
	x"63" when entrada = x"ee" else
	x"6d" when entrada = x"ef" else
	x"d7" when entrada = x"f0" else
	x"d9" when entrada = x"f1" else
	x"cb" when entrada = x"f2" else
	x"c5" when entrada = x"f3" else
	x"ef" when entrada = x"f4" else
	x"e1" when entrada = x"f5" else
	x"f3" when entrada = x"f6" else
	x"fd" when entrada = x"f7" else
	x"a7" when entrada = x"f8" else
	x"a9" when entrada = x"f9" else
	x"bb" when entrada = x"fa" else
	x"b5" when entrada = x"fb" else
	x"9f" when entrada = x"fc" else
	x"91" when entrada = x"fd" else
	x"83" when entrada = x"fe" else
	x"8d" when entrada = x"ff";
end catorze;
